module canvas


type SVGMatrix=[]f64
type Number =f64
type CanvasImageSource=string
type Point2D=[]f64
type Path2D=[]Point2D
type ImageDataSettings=map[string]string
type ImageData=string

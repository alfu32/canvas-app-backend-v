module utils

fn test_toast(){
	println(toast("you're toast !"))
}

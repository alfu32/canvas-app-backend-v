module geometry

pub struct TechnoLang{
	technoid string
	langid string
}
pub fn new_technolang() TechnoLang {
	return TechnoLang{}
}

module geometry

pub struct TechnoLang{
	technoid string
	langid string
}

module users

pub struct User{
	id string
	given_name string
	email string
	picture string
}


